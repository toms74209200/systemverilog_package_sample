/*=============================================================================
 * Title        : Package sample
 *
 * File Name    : foo_pkg.sv
 * Project      : 
 * Block        : 
 * Tree         : 
 * Designer     : toms74209200 <https://github.com/toms74209200>
 * Created      : 2020/01/09
 * License      : MIT License.
                  http://opensource.org/licenses/mit-license.php
 *============================================================================*/

package foo_pkg;

string str = "Hello, World!";

endpackage

import foo_pkg::*;